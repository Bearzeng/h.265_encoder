//-------------------------------------------------------------------
//
//  COPYRIGHT (C) 2014, VIPcore Group, Fudan University
//
//  THIS FILE MAY NOT BE MODIFIED OR REDISTRIBUTED WITHOUT THE
//  EXPRESSED WRITTEN CONSENT OF VIPcore Group
//
//  VIPcore       : http://soc.fudan.edu.cn/vip
//  IP Owner      : Yibo FAN
//  Contact       : fanyibo@fudan.edu.cn
//
//-------------------------------------------------------------------
//
//  Filename      : ime_systolic_array.v
//  Author        : Huang Lei Lei
//  Created       : 2014-12-10
//  Description   : systolic_array for reference and original pixels
//
//-------------------------------------------------------------------
//
//  Modification  : 2014-12-15
//  Description   : format of the input is merged
//                  order of the input is reversed (pixel_00_o should output the lastest input data)
//
//-------------------------------------------------------------------

`include "enc_defines.v"

module ime_systolic_array (
  // global
  clk             ,
  rstn            ,

  // shift_i
  shift_en_i      ,
  shift_data_i    ,

  // data_o
  pixel_00_o      ,
  pixel_01_o      ,
  pixel_02_o      ,
  pixel_03_o      ,
  pixel_04_o      ,
  pixel_05_o      ,
  pixel_06_o      ,
  pixel_07_o      ,
  pixel_08_o      ,
  pixel_09_o      ,
  pixel_10_o      ,
  pixel_11_o      ,
  pixel_12_o      ,
  pixel_13_o      ,
  pixel_14_o      ,
  pixel_15_o

/*  // pixel_00-03_00-63_o
  pixel_00_00_o    , pixel_01_00_o    , pixel_02_00_o    , pixel_03_00_o    ,
  pixel_00_01_o    , pixel_01_01_o    , pixel_02_01_o    , pixel_03_01_o    ,
  pixel_00_02_o    , pixel_01_02_o    , pixel_02_02_o    , pixel_03_02_o    ,
  pixel_00_03_o    , pixel_01_03_o    , pixel_02_03_o    , pixel_03_03_o    ,
  pixel_00_04_o    , pixel_01_04_o    , pixel_02_04_o    , pixel_03_04_o    ,
  pixel_00_05_o    , pixel_01_05_o    , pixel_02_05_o    , pixel_03_05_o    ,
  pixel_00_06_o    , pixel_01_06_o    , pixel_02_06_o    , pixel_03_06_o    ,
  pixel_00_07_o    , pixel_01_07_o    , pixel_02_07_o    , pixel_03_07_o    ,
  pixel_00_08_o    , pixel_01_08_o    , pixel_02_08_o    , pixel_03_08_o    ,
  pixel_00_09_o    , pixel_01_09_o    , pixel_02_09_o    , pixel_03_09_o    ,

  pixel_00_10_o    , pixel_01_10_o    , pixel_02_10_o    , pixel_03_10_o    ,
  pixel_00_11_o    , pixel_01_11_o    , pixel_02_11_o    , pixel_03_11_o    ,
  pixel_00_12_o    , pixel_01_12_o    , pixel_02_12_o    , pixel_03_12_o    ,
  pixel_00_13_o    , pixel_01_13_o    , pixel_02_13_o    , pixel_03_13_o    ,
  pixel_00_14_o    , pixel_01_14_o    , pixel_02_14_o    , pixel_03_14_o    ,
  pixel_00_15_o    , pixel_01_15_o    , pixel_02_15_o    , pixel_03_15_o    ,
  pixel_00_16_o    , pixel_01_16_o    , pixel_02_16_o    , pixel_03_16_o    ,
  pixel_00_17_o    , pixel_01_17_o    , pixel_02_17_o    , pixel_03_17_o    ,
  pixel_00_18_o    , pixel_01_18_o    , pixel_02_18_o    , pixel_03_18_o    ,
  pixel_00_19_o    , pixel_01_19_o    , pixel_02_19_o    , pixel_03_19_o    ,

  pixel_00_20_o    , pixel_01_20_o    , pixel_02_20_o    , pixel_03_20_o    ,
  pixel_00_21_o    , pixel_01_21_o    , pixel_02_21_o    , pixel_03_21_o    ,
  pixel_00_22_o    , pixel_01_22_o    , pixel_02_22_o    , pixel_03_22_o    ,
  pixel_00_23_o    , pixel_01_23_o    , pixel_02_23_o    , pixel_03_23_o    ,
  pixel_00_24_o    , pixel_01_24_o    , pixel_02_24_o    , pixel_03_24_o    ,
  pixel_00_25_o    , pixel_01_25_o    , pixel_02_25_o    , pixel_03_25_o    ,
  pixel_00_26_o    , pixel_01_26_o    , pixel_02_26_o    , pixel_03_26_o    ,
  pixel_00_27_o    , pixel_01_27_o    , pixel_02_27_o    , pixel_03_27_o    ,
  pixel_00_28_o    , pixel_01_28_o    , pixel_02_28_o    , pixel_03_28_o    ,
  pixel_00_29_o    , pixel_01_29_o    , pixel_02_29_o    , pixel_03_29_o    ,

  pixel_00_30_o    , pixel_01_30_o    , pixel_02_30_o    , pixel_03_30_o    ,
  pixel_00_31_o    , pixel_01_31_o    , pixel_02_31_o    , pixel_03_31_o    ,
  pixel_00_32_o    , pixel_01_32_o    , pixel_02_32_o    , pixel_03_32_o    ,
  pixel_00_33_o    , pixel_01_33_o    , pixel_02_33_o    , pixel_03_33_o    ,
  pixel_00_34_o    , pixel_01_34_o    , pixel_02_34_o    , pixel_03_34_o    ,
  pixel_00_35_o    , pixel_01_35_o    , pixel_02_35_o    , pixel_03_35_o    ,
  pixel_00_36_o    , pixel_01_36_o    , pixel_02_36_o    , pixel_03_36_o    ,
  pixel_00_37_o    , pixel_01_37_o    , pixel_02_37_o    , pixel_03_37_o    ,
  pixel_00_38_o    , pixel_01_38_o    , pixel_02_38_o    , pixel_03_38_o    ,
  pixel_00_39_o    , pixel_01_39_o    , pixel_02_39_o    , pixel_03_39_o    ,

  pixel_00_40_o    , pixel_01_40_o    , pixel_02_40_o    , pixel_03_40_o    ,
  pixel_00_41_o    , pixel_01_41_o    , pixel_02_41_o    , pixel_03_41_o    ,
  pixel_00_42_o    , pixel_01_42_o    , pixel_02_42_o    , pixel_03_42_o    ,
  pixel_00_43_o    , pixel_01_43_o    , pixel_02_43_o    , pixel_03_43_o    ,
  pixel_00_44_o    , pixel_01_44_o    , pixel_02_44_o    , pixel_03_44_o    ,
  pixel_00_45_o    , pixel_01_45_o    , pixel_02_45_o    , pixel_03_45_o    ,
  pixel_00_46_o    , pixel_01_46_o    , pixel_02_46_o    , pixel_03_46_o    ,
  pixel_00_47_o    , pixel_01_47_o    , pixel_02_47_o    , pixel_03_47_o    ,
  pixel_00_48_o    , pixel_01_48_o    , pixel_02_48_o    , pixel_03_48_o    ,
  pixel_00_49_o    , pixel_01_49_o    , pixel_02_49_o    , pixel_03_49_o    ,

  pixel_00_50_o    , pixel_01_50_o    , pixel_02_50_o    , pixel_03_50_o    ,
  pixel_00_51_o    , pixel_01_51_o    , pixel_02_51_o    , pixel_03_51_o    ,
  pixel_00_52_o    , pixel_01_52_o    , pixel_02_52_o    , pixel_03_52_o    ,
  pixel_00_53_o    , pixel_01_53_o    , pixel_02_53_o    , pixel_03_53_o    ,
  pixel_00_54_o    , pixel_01_54_o    , pixel_02_54_o    , pixel_03_54_o    ,
  pixel_00_55_o    , pixel_01_55_o    , pixel_02_55_o    , pixel_03_55_o    ,
  pixel_00_56_o    , pixel_01_56_o    , pixel_02_56_o    , pixel_03_56_o    ,
  pixel_00_57_o    , pixel_01_57_o    , pixel_02_57_o    , pixel_03_57_o    ,
  pixel_00_58_o    , pixel_01_58_o    , pixel_02_58_o    , pixel_03_58_o    ,
  pixel_00_59_o    , pixel_01_59_o    , pixel_02_59_o    , pixel_03_59_o    ,

  pixel_00_60_o    , pixel_01_60_o    , pixel_02_60_o    , pixel_03_60_o    ,
  pixel_00_61_o    , pixel_01_61_o    , pixel_02_61_o    , pixel_03_61_o    ,
  pixel_00_62_o    , pixel_01_62_o    , pixel_02_62_o    , pixel_03_62_o    ,
  pixel_00_63_o    , pixel_01_63_o    , pixel_02_63_o    , pixel_03_63_o    ,

  // pixel_04-07_00-63_o
  pixel_04_00_o    , pixel_05_00_o    , pixel_06_00_o    , pixel_07_00_o    ,
  pixel_04_01_o    , pixel_05_01_o    , pixel_06_01_o    , pixel_07_01_o    ,
  pixel_04_02_o    , pixel_05_02_o    , pixel_06_02_o    , pixel_07_02_o    ,
  pixel_04_03_o    , pixel_05_03_o    , pixel_06_03_o    , pixel_07_03_o    ,
  pixel_04_04_o    , pixel_05_04_o    , pixel_06_04_o    , pixel_07_04_o    ,
  pixel_04_05_o    , pixel_05_05_o    , pixel_06_05_o    , pixel_07_05_o    ,
  pixel_04_06_o    , pixel_05_06_o    , pixel_06_06_o    , pixel_07_06_o    ,
  pixel_04_07_o    , pixel_05_07_o    , pixel_06_07_o    , pixel_07_07_o    ,
  pixel_04_08_o    , pixel_05_08_o    , pixel_06_08_o    , pixel_07_08_o    ,
  pixel_04_09_o    , pixel_05_09_o    , pixel_06_09_o    , pixel_07_09_o    ,

  pixel_04_10_o    , pixel_05_10_o    , pixel_06_10_o    , pixel_07_10_o    ,
  pixel_04_11_o    , pixel_05_11_o    , pixel_06_11_o    , pixel_07_11_o    ,
  pixel_04_12_o    , pixel_05_12_o    , pixel_06_12_o    , pixel_07_12_o    ,
  pixel_04_13_o    , pixel_05_13_o    , pixel_06_13_o    , pixel_07_13_o    ,
  pixel_04_14_o    , pixel_05_14_o    , pixel_06_14_o    , pixel_07_14_o    ,
  pixel_04_15_o    , pixel_05_15_o    , pixel_06_15_o    , pixel_07_15_o    ,
  pixel_04_16_o    , pixel_05_16_o    , pixel_06_16_o    , pixel_07_16_o    ,
  pixel_04_17_o    , pixel_05_17_o    , pixel_06_17_o    , pixel_07_17_o    ,
  pixel_04_18_o    , pixel_05_18_o    , pixel_06_18_o    , pixel_07_18_o    ,
  pixel_04_19_o    , pixel_05_19_o    , pixel_06_19_o    , pixel_07_19_o    ,

  pixel_04_20_o    , pixel_05_20_o    , pixel_06_20_o    , pixel_07_20_o    ,
  pixel_04_21_o    , pixel_05_21_o    , pixel_06_21_o    , pixel_07_21_o    ,
  pixel_04_22_o    , pixel_05_22_o    , pixel_06_22_o    , pixel_07_22_o    ,
  pixel_04_23_o    , pixel_05_23_o    , pixel_06_23_o    , pixel_07_23_o    ,
  pixel_04_24_o    , pixel_05_24_o    , pixel_06_24_o    , pixel_07_24_o    ,
  pixel_04_25_o    , pixel_05_25_o    , pixel_06_25_o    , pixel_07_25_o    ,
  pixel_04_26_o    , pixel_05_26_o    , pixel_06_26_o    , pixel_07_26_o    ,
  pixel_04_27_o    , pixel_05_27_o    , pixel_06_27_o    , pixel_07_27_o    ,
  pixel_04_28_o    , pixel_05_28_o    , pixel_06_28_o    , pixel_07_28_o    ,
  pixel_04_29_o    , pixel_05_29_o    , pixel_06_29_o    , pixel_07_29_o    ,

  pixel_04_30_o    , pixel_05_30_o    , pixel_06_30_o    , pixel_07_30_o    ,
  pixel_04_31_o    , pixel_05_31_o    , pixel_06_31_o    , pixel_07_31_o    ,
  pixel_04_32_o    , pixel_05_32_o    , pixel_06_32_o    , pixel_07_32_o    ,
  pixel_04_33_o    , pixel_05_33_o    , pixel_06_33_o    , pixel_07_33_o    ,
  pixel_04_34_o    , pixel_05_34_o    , pixel_06_34_o    , pixel_07_34_o    ,
  pixel_04_35_o    , pixel_05_35_o    , pixel_06_35_o    , pixel_07_35_o    ,
  pixel_04_36_o    , pixel_05_36_o    , pixel_06_36_o    , pixel_07_36_o    ,
  pixel_04_37_o    , pixel_05_37_o    , pixel_06_37_o    , pixel_07_37_o    ,
  pixel_04_38_o    , pixel_05_38_o    , pixel_06_38_o    , pixel_07_38_o    ,
  pixel_04_39_o    , pixel_05_39_o    , pixel_06_39_o    , pixel_07_39_o    ,

  pixel_04_40_o    , pixel_05_40_o    , pixel_06_40_o    , pixel_07_40_o    ,
  pixel_04_41_o    , pixel_05_41_o    , pixel_06_41_o    , pixel_07_41_o    ,
  pixel_04_42_o    , pixel_05_42_o    , pixel_06_42_o    , pixel_07_42_o    ,
  pixel_04_43_o    , pixel_05_43_o    , pixel_06_43_o    , pixel_07_43_o    ,
  pixel_04_44_o    , pixel_05_44_o    , pixel_06_44_o    , pixel_07_44_o    ,
  pixel_04_45_o    , pixel_05_45_o    , pixel_06_45_o    , pixel_07_45_o    ,
  pixel_04_46_o    , pixel_05_46_o    , pixel_06_46_o    , pixel_07_46_o    ,
  pixel_04_47_o    , pixel_05_47_o    , pixel_06_47_o    , pixel_07_47_o    ,
  pixel_04_48_o    , pixel_05_48_o    , pixel_06_48_o    , pixel_07_48_o    ,
  pixel_04_49_o    , pixel_05_49_o    , pixel_06_49_o    , pixel_07_49_o    ,

  pixel_04_50_o    , pixel_05_50_o    , pixel_06_50_o    , pixel_07_50_o    ,
  pixel_04_51_o    , pixel_05_51_o    , pixel_06_51_o    , pixel_07_51_o    ,
  pixel_04_52_o    , pixel_05_52_o    , pixel_06_52_o    , pixel_07_52_o    ,
  pixel_04_53_o    , pixel_05_53_o    , pixel_06_53_o    , pixel_07_53_o    ,
  pixel_04_54_o    , pixel_05_54_o    , pixel_06_54_o    , pixel_07_54_o    ,
  pixel_04_55_o    , pixel_05_55_o    , pixel_06_55_o    , pixel_07_55_o    ,
  pixel_04_56_o    , pixel_05_56_o    , pixel_06_56_o    , pixel_07_56_o    ,
  pixel_04_57_o    , pixel_05_57_o    , pixel_06_57_o    , pixel_07_57_o    ,
  pixel_04_58_o    , pixel_05_58_o    , pixel_06_58_o    , pixel_07_58_o    ,
  pixel_04_59_o    , pixel_05_59_o    , pixel_06_59_o    , pixel_07_59_o    ,

  pixel_04_60_o    , pixel_05_60_o    , pixel_06_60_o    , pixel_07_60_o    ,
  pixel_04_61_o    , pixel_05_61_o    , pixel_06_61_o    , pixel_07_61_o    ,
  pixel_04_62_o    , pixel_05_62_o    , pixel_06_62_o    , pixel_07_62_o    ,
  pixel_04_63_o    , pixel_05_63_o    , pixel_06_63_o    , pixel_07_63_o    ,

  // pixel_08-11_00-63_o
  pixel_08_00_o    , pixel_09_00_o    , pixel_10_00_o    , pixel_11_00_o    ,
  pixel_08_01_o    , pixel_09_01_o    , pixel_10_01_o    , pixel_11_01_o    ,
  pixel_08_02_o    , pixel_09_02_o    , pixel_10_02_o    , pixel_11_02_o    ,
  pixel_08_03_o    , pixel_09_03_o    , pixel_10_03_o    , pixel_11_03_o    ,
  pixel_08_04_o    , pixel_09_04_o    , pixel_10_04_o    , pixel_11_04_o    ,
  pixel_08_05_o    , pixel_09_05_o    , pixel_10_05_o    , pixel_11_05_o    ,
  pixel_08_06_o    , pixel_09_06_o    , pixel_10_06_o    , pixel_11_06_o    ,
  pixel_08_07_o    , pixel_09_07_o    , pixel_10_07_o    , pixel_11_07_o    ,
  pixel_08_08_o    , pixel_09_08_o    , pixel_10_08_o    , pixel_11_08_o    ,
  pixel_08_09_o    , pixel_09_09_o    , pixel_10_09_o    , pixel_11_09_o    ,

  pixel_08_10_o    , pixel_09_10_o    , pixel_10_10_o    , pixel_11_10_o    ,
  pixel_08_11_o    , pixel_09_11_o    , pixel_10_11_o    , pixel_11_11_o    ,
  pixel_08_12_o    , pixel_09_12_o    , pixel_10_12_o    , pixel_11_12_o    ,
  pixel_08_13_o    , pixel_09_13_o    , pixel_10_13_o    , pixel_11_13_o    ,
  pixel_08_14_o    , pixel_09_14_o    , pixel_10_14_o    , pixel_11_14_o    ,
  pixel_08_15_o    , pixel_09_15_o    , pixel_10_15_o    , pixel_11_15_o    ,
  pixel_08_16_o    , pixel_09_16_o    , pixel_10_16_o    , pixel_11_16_o    ,
  pixel_08_17_o    , pixel_09_17_o    , pixel_10_17_o    , pixel_11_17_o    ,
  pixel_08_18_o    , pixel_09_18_o    , pixel_10_18_o    , pixel_11_18_o    ,
  pixel_08_19_o    , pixel_09_19_o    , pixel_10_19_o    , pixel_11_19_o    ,

  pixel_08_20_o    , pixel_09_20_o    , pixel_10_20_o    , pixel_11_20_o    ,
  pixel_08_21_o    , pixel_09_21_o    , pixel_10_21_o    , pixel_11_21_o    ,
  pixel_08_22_o    , pixel_09_22_o    , pixel_10_22_o    , pixel_11_22_o    ,
  pixel_08_23_o    , pixel_09_23_o    , pixel_10_23_o    , pixel_11_23_o    ,
  pixel_08_24_o    , pixel_09_24_o    , pixel_10_24_o    , pixel_11_24_o    ,
  pixel_08_25_o    , pixel_09_25_o    , pixel_10_25_o    , pixel_11_25_o    ,
  pixel_08_26_o    , pixel_09_26_o    , pixel_10_26_o    , pixel_11_26_o    ,
  pixel_08_27_o    , pixel_09_27_o    , pixel_10_27_o    , pixel_11_27_o    ,
  pixel_08_28_o    , pixel_09_28_o    , pixel_10_28_o    , pixel_11_28_o    ,
  pixel_08_29_o    , pixel_09_29_o    , pixel_10_29_o    , pixel_11_29_o    ,

  pixel_08_30_o    , pixel_09_30_o    , pixel_10_30_o    , pixel_11_30_o    ,
  pixel_08_31_o    , pixel_09_31_o    , pixel_10_31_o    , pixel_11_31_o    ,
  pixel_08_32_o    , pixel_09_32_o    , pixel_10_32_o    , pixel_11_32_o    ,
  pixel_08_33_o    , pixel_09_33_o    , pixel_10_33_o    , pixel_11_33_o    ,
  pixel_08_34_o    , pixel_09_34_o    , pixel_10_34_o    , pixel_11_34_o    ,
  pixel_08_35_o    , pixel_09_35_o    , pixel_10_35_o    , pixel_11_35_o    ,
  pixel_08_36_o    , pixel_09_36_o    , pixel_10_36_o    , pixel_11_36_o    ,
  pixel_08_37_o    , pixel_09_37_o    , pixel_10_37_o    , pixel_11_37_o    ,
  pixel_08_38_o    , pixel_09_38_o    , pixel_10_38_o    , pixel_11_38_o    ,
  pixel_08_39_o    , pixel_09_39_o    , pixel_10_39_o    , pixel_11_39_o    ,

  pixel_08_40_o    , pixel_09_40_o    , pixel_10_40_o    , pixel_11_40_o    ,
  pixel_08_41_o    , pixel_09_41_o    , pixel_10_41_o    , pixel_11_41_o    ,
  pixel_08_42_o    , pixel_09_42_o    , pixel_10_42_o    , pixel_11_42_o    ,
  pixel_08_43_o    , pixel_09_43_o    , pixel_10_43_o    , pixel_11_43_o    ,
  pixel_08_44_o    , pixel_09_44_o    , pixel_10_44_o    , pixel_11_44_o    ,
  pixel_08_45_o    , pixel_09_45_o    , pixel_10_45_o    , pixel_11_45_o    ,
  pixel_08_46_o    , pixel_09_46_o    , pixel_10_46_o    , pixel_11_46_o    ,
  pixel_08_47_o    , pixel_09_47_o    , pixel_10_47_o    , pixel_11_47_o    ,
  pixel_08_48_o    , pixel_09_48_o    , pixel_10_48_o    , pixel_11_48_o    ,
  pixel_08_49_o    , pixel_09_49_o    , pixel_10_49_o    , pixel_11_49_o    ,

  pixel_08_50_o    , pixel_09_50_o    , pixel_10_50_o    , pixel_11_50_o    ,
  pixel_08_51_o    , pixel_09_51_o    , pixel_10_51_o    , pixel_11_51_o    ,
  pixel_08_52_o    , pixel_09_52_o    , pixel_10_52_o    , pixel_11_52_o    ,
  pixel_08_53_o    , pixel_09_53_o    , pixel_10_53_o    , pixel_11_53_o    ,
  pixel_08_54_o    , pixel_09_54_o    , pixel_10_54_o    , pixel_11_54_o    ,
  pixel_08_55_o    , pixel_09_55_o    , pixel_10_55_o    , pixel_11_55_o    ,
  pixel_08_56_o    , pixel_09_56_o    , pixel_10_56_o    , pixel_11_56_o    ,
  pixel_08_57_o    , pixel_09_57_o    , pixel_10_57_o    , pixel_11_57_o    ,
  pixel_08_58_o    , pixel_09_58_o    , pixel_10_58_o    , pixel_11_58_o    ,
  pixel_08_59_o    , pixel_09_59_o    , pixel_10_59_o    , pixel_11_59_o    ,

  pixel_08_60_o    , pixel_09_60_o    , pixel_10_60_o    , pixel_11_60_o    ,
  pixel_08_61_o    , pixel_09_61_o    , pixel_10_61_o    , pixel_11_61_o    ,
  pixel_08_62_o    , pixel_09_62_o    , pixel_10_62_o    , pixel_11_62_o    ,
  pixel_08_63_o    , pixel_09_63_o    , pixel_10_63_o    , pixel_11_63_o    ,

  // pixel_12-15_00-63_o
  pixel_12_00_o    , pixel_13_00_o    , pixel_14_00_o    , pixel_15_00_o    ,
  pixel_12_01_o    , pixel_13_01_o    , pixel_14_01_o    , pixel_15_01_o    ,
  pixel_12_02_o    , pixel_13_02_o    , pixel_14_02_o    , pixel_15_02_o    ,
  pixel_12_03_o    , pixel_13_03_o    , pixel_14_03_o    , pixel_15_03_o    ,
  pixel_12_04_o    , pixel_13_04_o    , pixel_14_04_o    , pixel_15_04_o    ,
  pixel_12_05_o    , pixel_13_05_o    , pixel_14_05_o    , pixel_15_05_o    ,
  pixel_12_06_o    , pixel_13_06_o    , pixel_14_06_o    , pixel_15_06_o    ,
  pixel_12_07_o    , pixel_13_07_o    , pixel_14_07_o    , pixel_15_07_o    ,
  pixel_12_08_o    , pixel_13_08_o    , pixel_14_08_o    , pixel_15_08_o    ,
  pixel_12_09_o    , pixel_13_09_o    , pixel_14_09_o    , pixel_15_09_o    ,

  pixel_12_10_o    , pixel_13_10_o    , pixel_14_10_o    , pixel_15_10_o    ,
  pixel_12_11_o    , pixel_13_11_o    , pixel_14_11_o    , pixel_15_11_o    ,
  pixel_12_12_o    , pixel_13_12_o    , pixel_14_12_o    , pixel_15_12_o    ,
  pixel_12_13_o    , pixel_13_13_o    , pixel_14_13_o    , pixel_15_13_o    ,
  pixel_12_14_o    , pixel_13_14_o    , pixel_14_14_o    , pixel_15_14_o    ,
  pixel_12_15_o    , pixel_13_15_o    , pixel_14_15_o    , pixel_15_15_o    ,
  pixel_12_16_o    , pixel_13_16_o    , pixel_14_16_o    , pixel_15_16_o    ,
  pixel_12_17_o    , pixel_13_17_o    , pixel_14_17_o    , pixel_15_17_o    ,
  pixel_12_18_o    , pixel_13_18_o    , pixel_14_18_o    , pixel_15_18_o    ,
  pixel_12_19_o    , pixel_13_19_o    , pixel_14_19_o    , pixel_15_19_o    ,

  pixel_12_20_o    , pixel_13_20_o    , pixel_14_20_o    , pixel_15_20_o    ,
  pixel_12_21_o    , pixel_13_21_o    , pixel_14_21_o    , pixel_15_21_o    ,
  pixel_12_22_o    , pixel_13_22_o    , pixel_14_22_o    , pixel_15_22_o    ,
  pixel_12_23_o    , pixel_13_23_o    , pixel_14_23_o    , pixel_15_23_o    ,
  pixel_12_24_o    , pixel_13_24_o    , pixel_14_24_o    , pixel_15_24_o    ,
  pixel_12_25_o    , pixel_13_25_o    , pixel_14_25_o    , pixel_15_25_o    ,
  pixel_12_26_o    , pixel_13_26_o    , pixel_14_26_o    , pixel_15_26_o    ,
  pixel_12_27_o    , pixel_13_27_o    , pixel_14_27_o    , pixel_15_27_o    ,
  pixel_12_28_o    , pixel_13_28_o    , pixel_14_28_o    , pixel_15_28_o    ,
  pixel_12_29_o    , pixel_13_29_o    , pixel_14_29_o    , pixel_15_29_o    ,

  pixel_12_30_o    , pixel_13_30_o    , pixel_14_30_o    , pixel_15_30_o    ,
  pixel_12_31_o    , pixel_13_31_o    , pixel_14_31_o    , pixel_15_31_o    ,
  pixel_12_32_o    , pixel_13_32_o    , pixel_14_32_o    , pixel_15_32_o    ,
  pixel_12_33_o    , pixel_13_33_o    , pixel_14_33_o    , pixel_15_33_o    ,
  pixel_12_34_o    , pixel_13_34_o    , pixel_14_34_o    , pixel_15_34_o    ,
  pixel_12_35_o    , pixel_13_35_o    , pixel_14_35_o    , pixel_15_35_o    ,
  pixel_12_36_o    , pixel_13_36_o    , pixel_14_36_o    , pixel_15_36_o    ,
  pixel_12_37_o    , pixel_13_37_o    , pixel_14_37_o    , pixel_15_37_o    ,
  pixel_12_38_o    , pixel_13_38_o    , pixel_14_38_o    , pixel_15_38_o    ,
  pixel_12_39_o    , pixel_13_39_o    , pixel_14_39_o    , pixel_15_39_o    ,

  pixel_12_40_o    , pixel_13_40_o    , pixel_14_40_o    , pixel_15_40_o    ,
  pixel_12_41_o    , pixel_13_41_o    , pixel_14_41_o    , pixel_15_41_o    ,
  pixel_12_42_o    , pixel_13_42_o    , pixel_14_42_o    , pixel_15_42_o    ,
  pixel_12_43_o    , pixel_13_43_o    , pixel_14_43_o    , pixel_15_43_o    ,
  pixel_12_44_o    , pixel_13_44_o    , pixel_14_44_o    , pixel_15_44_o    ,
  pixel_12_45_o    , pixel_13_45_o    , pixel_14_45_o    , pixel_15_45_o    ,
  pixel_12_46_o    , pixel_13_46_o    , pixel_14_46_o    , pixel_15_46_o    ,
  pixel_12_47_o    , pixel_13_47_o    , pixel_14_47_o    , pixel_15_47_o    ,
  pixel_12_48_o    , pixel_13_48_o    , pixel_14_48_o    , pixel_15_48_o    ,
  pixel_12_49_o    , pixel_13_49_o    , pixel_14_49_o    , pixel_15_49_o    ,

  pixel_12_50_o    , pixel_13_50_o    , pixel_14_50_o    , pixel_15_50_o    ,
  pixel_12_51_o    , pixel_13_51_o    , pixel_14_51_o    , pixel_15_51_o    ,
  pixel_12_52_o    , pixel_13_52_o    , pixel_14_52_o    , pixel_15_52_o    ,
  pixel_12_53_o    , pixel_13_53_o    , pixel_14_53_o    , pixel_15_53_o    ,
  pixel_12_54_o    , pixel_13_54_o    , pixel_14_54_o    , pixel_15_54_o    ,
  pixel_12_55_o    , pixel_13_55_o    , pixel_14_55_o    , pixel_15_55_o    ,
  pixel_12_56_o    , pixel_13_56_o    , pixel_14_56_o    , pixel_15_56_o    ,
  pixel_12_57_o    , pixel_13_57_o    , pixel_14_57_o    , pixel_15_57_o    ,
  pixel_12_58_o    , pixel_13_58_o    , pixel_14_58_o    , pixel_15_58_o    ,
  pixel_12_59_o    , pixel_13_59_o    , pixel_14_59_o    , pixel_15_59_o    ,

  pixel_12_60_o    , pixel_13_60_o    , pixel_14_60_o    , pixel_15_60_o    ,
  pixel_12_61_o    , pixel_13_61_o    , pixel_14_61_o    , pixel_15_61_o    ,
  pixel_12_62_o    , pixel_13_62_o    , pixel_14_62_o    , pixel_15_62_o    ,
  pixel_12_63_o    , pixel_13_63_o    , pixel_14_63_o    , pixel_15_63_o
*/  );


//*** PARAMETER DECLARATION ****************************************************


//*** INPUT/OUTPUT DECLARATION *************************************************

  // global
  input                             clk             ;
  input                             rstn            ;

  // shift_i
  input                             shift_en_i      ;
  input  [`PIXEL_WIDTH*64-1 : 0]    shift_data_i    ;

  // data_o
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_00_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_01_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_02_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_03_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_04_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_05_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_06_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_07_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_08_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_09_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_10_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_11_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_12_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_13_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_14_o      ;
  output [`PIXEL_WIDTH*64-1 : 0]    pixel_15_o      ;

/*  // pixel_00-03_00-63_o
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_00_o    , pixel_01_00_o    , pixel_02_00_o    , pixel_03_00_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_01_o    , pixel_01_01_o    , pixel_02_01_o    , pixel_03_01_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_02_o    , pixel_01_02_o    , pixel_02_02_o    , pixel_03_02_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_03_o    , pixel_01_03_o    , pixel_02_03_o    , pixel_03_03_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_04_o    , pixel_01_04_o    , pixel_02_04_o    , pixel_03_04_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_05_o    , pixel_01_05_o    , pixel_02_05_o    , pixel_03_05_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_06_o    , pixel_01_06_o    , pixel_02_06_o    , pixel_03_06_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_07_o    , pixel_01_07_o    , pixel_02_07_o    , pixel_03_07_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_08_o    , pixel_01_08_o    , pixel_02_08_o    , pixel_03_08_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_09_o    , pixel_01_09_o    , pixel_02_09_o    , pixel_03_09_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_00_10_o    , pixel_01_10_o    , pixel_02_10_o    , pixel_03_10_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_11_o    , pixel_01_11_o    , pixel_02_11_o    , pixel_03_11_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_12_o    , pixel_01_12_o    , pixel_02_12_o    , pixel_03_12_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_13_o    , pixel_01_13_o    , pixel_02_13_o    , pixel_03_13_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_14_o    , pixel_01_14_o    , pixel_02_14_o    , pixel_03_14_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_15_o    , pixel_01_15_o    , pixel_02_15_o    , pixel_03_15_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_16_o    , pixel_01_16_o    , pixel_02_16_o    , pixel_03_16_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_17_o    , pixel_01_17_o    , pixel_02_17_o    , pixel_03_17_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_18_o    , pixel_01_18_o    , pixel_02_18_o    , pixel_03_18_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_19_o    , pixel_01_19_o    , pixel_02_19_o    , pixel_03_19_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_00_20_o    , pixel_01_20_o    , pixel_02_20_o    , pixel_03_20_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_21_o    , pixel_01_21_o    , pixel_02_21_o    , pixel_03_21_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_22_o    , pixel_01_22_o    , pixel_02_22_o    , pixel_03_22_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_23_o    , pixel_01_23_o    , pixel_02_23_o    , pixel_03_23_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_24_o    , pixel_01_24_o    , pixel_02_24_o    , pixel_03_24_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_25_o    , pixel_01_25_o    , pixel_02_25_o    , pixel_03_25_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_26_o    , pixel_01_26_o    , pixel_02_26_o    , pixel_03_26_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_27_o    , pixel_01_27_o    , pixel_02_27_o    , pixel_03_27_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_28_o    , pixel_01_28_o    , pixel_02_28_o    , pixel_03_28_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_29_o    , pixel_01_29_o    , pixel_02_29_o    , pixel_03_29_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_00_30_o    , pixel_01_30_o    , pixel_02_30_o    , pixel_03_30_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_31_o    , pixel_01_31_o    , pixel_02_31_o    , pixel_03_31_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_32_o    , pixel_01_32_o    , pixel_02_32_o    , pixel_03_32_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_33_o    , pixel_01_33_o    , pixel_02_33_o    , pixel_03_33_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_34_o    , pixel_01_34_o    , pixel_02_34_o    , pixel_03_34_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_35_o    , pixel_01_35_o    , pixel_02_35_o    , pixel_03_35_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_36_o    , pixel_01_36_o    , pixel_02_36_o    , pixel_03_36_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_37_o    , pixel_01_37_o    , pixel_02_37_o    , pixel_03_37_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_38_o    , pixel_01_38_o    , pixel_02_38_o    , pixel_03_38_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_39_o    , pixel_01_39_o    , pixel_02_39_o    , pixel_03_39_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_00_40_o    , pixel_01_40_o    , pixel_02_40_o    , pixel_03_40_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_41_o    , pixel_01_41_o    , pixel_02_41_o    , pixel_03_41_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_42_o    , pixel_01_42_o    , pixel_02_42_o    , pixel_03_42_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_43_o    , pixel_01_43_o    , pixel_02_43_o    , pixel_03_43_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_44_o    , pixel_01_44_o    , pixel_02_44_o    , pixel_03_44_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_45_o    , pixel_01_45_o    , pixel_02_45_o    , pixel_03_45_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_46_o    , pixel_01_46_o    , pixel_02_46_o    , pixel_03_46_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_47_o    , pixel_01_47_o    , pixel_02_47_o    , pixel_03_47_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_48_o    , pixel_01_48_o    , pixel_02_48_o    , pixel_03_48_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_49_o    , pixel_01_49_o    , pixel_02_49_o    , pixel_03_49_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_00_50_o    , pixel_01_50_o    , pixel_02_50_o    , pixel_03_50_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_51_o    , pixel_01_51_o    , pixel_02_51_o    , pixel_03_51_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_52_o    , pixel_01_52_o    , pixel_02_52_o    , pixel_03_52_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_53_o    , pixel_01_53_o    , pixel_02_53_o    , pixel_03_53_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_54_o    , pixel_01_54_o    , pixel_02_54_o    , pixel_03_54_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_55_o    , pixel_01_55_o    , pixel_02_55_o    , pixel_03_55_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_56_o    , pixel_01_56_o    , pixel_02_56_o    , pixel_03_56_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_57_o    , pixel_01_57_o    , pixel_02_57_o    , pixel_03_57_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_58_o    , pixel_01_58_o    , pixel_02_58_o    , pixel_03_58_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_59_o    , pixel_01_59_o    , pixel_02_59_o    , pixel_03_59_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_00_60_o    , pixel_01_60_o    , pixel_02_60_o    , pixel_03_60_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_61_o    , pixel_01_61_o    , pixel_02_61_o    , pixel_03_61_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_62_o    , pixel_01_62_o    , pixel_02_62_o    , pixel_03_62_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_00_63_o    , pixel_01_63_o    , pixel_02_63_o    , pixel_03_63_o    ;

  // pixel_04-07_00-63_o
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_00_o    , pixel_05_00_o    , pixel_06_00_o    , pixel_07_00_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_01_o    , pixel_05_01_o    , pixel_06_01_o    , pixel_07_01_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_02_o    , pixel_05_02_o    , pixel_06_02_o    , pixel_07_02_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_03_o    , pixel_05_03_o    , pixel_06_03_o    , pixel_07_03_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_04_o    , pixel_05_04_o    , pixel_06_04_o    , pixel_07_04_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_05_o    , pixel_05_05_o    , pixel_06_05_o    , pixel_07_05_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_06_o    , pixel_05_06_o    , pixel_06_06_o    , pixel_07_06_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_07_o    , pixel_05_07_o    , pixel_06_07_o    , pixel_07_07_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_08_o    , pixel_05_08_o    , pixel_06_08_o    , pixel_07_08_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_09_o    , pixel_05_09_o    , pixel_06_09_o    , pixel_07_09_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_04_10_o    , pixel_05_10_o    , pixel_06_10_o    , pixel_07_10_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_11_o    , pixel_05_11_o    , pixel_06_11_o    , pixel_07_11_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_12_o    , pixel_05_12_o    , pixel_06_12_o    , pixel_07_12_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_13_o    , pixel_05_13_o    , pixel_06_13_o    , pixel_07_13_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_14_o    , pixel_05_14_o    , pixel_06_14_o    , pixel_07_14_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_15_o    , pixel_05_15_o    , pixel_06_15_o    , pixel_07_15_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_16_o    , pixel_05_16_o    , pixel_06_16_o    , pixel_07_16_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_17_o    , pixel_05_17_o    , pixel_06_17_o    , pixel_07_17_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_18_o    , pixel_05_18_o    , pixel_06_18_o    , pixel_07_18_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_19_o    , pixel_05_19_o    , pixel_06_19_o    , pixel_07_19_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_04_20_o    , pixel_05_20_o    , pixel_06_20_o    , pixel_07_20_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_21_o    , pixel_05_21_o    , pixel_06_21_o    , pixel_07_21_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_22_o    , pixel_05_22_o    , pixel_06_22_o    , pixel_07_22_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_23_o    , pixel_05_23_o    , pixel_06_23_o    , pixel_07_23_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_24_o    , pixel_05_24_o    , pixel_06_24_o    , pixel_07_24_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_25_o    , pixel_05_25_o    , pixel_06_25_o    , pixel_07_25_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_26_o    , pixel_05_26_o    , pixel_06_26_o    , pixel_07_26_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_27_o    , pixel_05_27_o    , pixel_06_27_o    , pixel_07_27_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_28_o    , pixel_05_28_o    , pixel_06_28_o    , pixel_07_28_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_29_o    , pixel_05_29_o    , pixel_06_29_o    , pixel_07_29_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_04_30_o    , pixel_05_30_o    , pixel_06_30_o    , pixel_07_30_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_31_o    , pixel_05_31_o    , pixel_06_31_o    , pixel_07_31_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_32_o    , pixel_05_32_o    , pixel_06_32_o    , pixel_07_32_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_33_o    , pixel_05_33_o    , pixel_06_33_o    , pixel_07_33_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_34_o    , pixel_05_34_o    , pixel_06_34_o    , pixel_07_34_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_35_o    , pixel_05_35_o    , pixel_06_35_o    , pixel_07_35_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_36_o    , pixel_05_36_o    , pixel_06_36_o    , pixel_07_36_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_37_o    , pixel_05_37_o    , pixel_06_37_o    , pixel_07_37_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_38_o    , pixel_05_38_o    , pixel_06_38_o    , pixel_07_38_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_39_o    , pixel_05_39_o    , pixel_06_39_o    , pixel_07_39_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_04_40_o    , pixel_05_40_o    , pixel_06_40_o    , pixel_07_40_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_41_o    , pixel_05_41_o    , pixel_06_41_o    , pixel_07_41_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_42_o    , pixel_05_42_o    , pixel_06_42_o    , pixel_07_42_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_43_o    , pixel_05_43_o    , pixel_06_43_o    , pixel_07_43_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_44_o    , pixel_05_44_o    , pixel_06_44_o    , pixel_07_44_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_45_o    , pixel_05_45_o    , pixel_06_45_o    , pixel_07_45_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_46_o    , pixel_05_46_o    , pixel_06_46_o    , pixel_07_46_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_47_o    , pixel_05_47_o    , pixel_06_47_o    , pixel_07_47_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_48_o    , pixel_05_48_o    , pixel_06_48_o    , pixel_07_48_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_49_o    , pixel_05_49_o    , pixel_06_49_o    , pixel_07_49_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_04_50_o    , pixel_05_50_o    , pixel_06_50_o    , pixel_07_50_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_51_o    , pixel_05_51_o    , pixel_06_51_o    , pixel_07_51_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_52_o    , pixel_05_52_o    , pixel_06_52_o    , pixel_07_52_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_53_o    , pixel_05_53_o    , pixel_06_53_o    , pixel_07_53_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_54_o    , pixel_05_54_o    , pixel_06_54_o    , pixel_07_54_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_55_o    , pixel_05_55_o    , pixel_06_55_o    , pixel_07_55_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_56_o    , pixel_05_56_o    , pixel_06_56_o    , pixel_07_56_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_57_o    , pixel_05_57_o    , pixel_06_57_o    , pixel_07_57_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_58_o    , pixel_05_58_o    , pixel_06_58_o    , pixel_07_58_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_59_o    , pixel_05_59_o    , pixel_06_59_o    , pixel_07_59_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_04_60_o    , pixel_05_60_o    , pixel_06_60_o    , pixel_07_60_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_61_o    , pixel_05_61_o    , pixel_06_61_o    , pixel_07_61_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_62_o    , pixel_05_62_o    , pixel_06_62_o    , pixel_07_62_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_04_63_o    , pixel_05_63_o    , pixel_06_63_o    , pixel_07_63_o    ;

  // pixel_08-11_00-63_o
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_00_o    , pixel_09_00_o    , pixel_10_00_o    , pixel_11_00_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_01_o    , pixel_09_01_o    , pixel_10_01_o    , pixel_11_01_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_02_o    , pixel_09_02_o    , pixel_10_02_o    , pixel_11_02_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_03_o    , pixel_09_03_o    , pixel_10_03_o    , pixel_11_03_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_04_o    , pixel_09_04_o    , pixel_10_04_o    , pixel_11_04_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_05_o    , pixel_09_05_o    , pixel_10_05_o    , pixel_11_05_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_06_o    , pixel_09_06_o    , pixel_10_06_o    , pixel_11_06_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_07_o    , pixel_09_07_o    , pixel_10_07_o    , pixel_11_07_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_08_o    , pixel_09_08_o    , pixel_10_08_o    , pixel_11_08_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_09_o    , pixel_09_09_o    , pixel_10_09_o    , pixel_11_09_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_08_10_o    , pixel_09_10_o    , pixel_10_10_o    , pixel_11_10_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_11_o    , pixel_09_11_o    , pixel_10_11_o    , pixel_11_11_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_12_o    , pixel_09_12_o    , pixel_10_12_o    , pixel_11_12_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_13_o    , pixel_09_13_o    , pixel_10_13_o    , pixel_11_13_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_14_o    , pixel_09_14_o    , pixel_10_14_o    , pixel_11_14_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_15_o    , pixel_09_15_o    , pixel_10_15_o    , pixel_11_15_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_16_o    , pixel_09_16_o    , pixel_10_16_o    , pixel_11_16_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_17_o    , pixel_09_17_o    , pixel_10_17_o    , pixel_11_17_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_18_o    , pixel_09_18_o    , pixel_10_18_o    , pixel_11_18_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_19_o    , pixel_09_19_o    , pixel_10_19_o    , pixel_11_19_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_08_20_o    , pixel_09_20_o    , pixel_10_20_o    , pixel_11_20_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_21_o    , pixel_09_21_o    , pixel_10_21_o    , pixel_11_21_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_22_o    , pixel_09_22_o    , pixel_10_22_o    , pixel_11_22_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_23_o    , pixel_09_23_o    , pixel_10_23_o    , pixel_11_23_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_24_o    , pixel_09_24_o    , pixel_10_24_o    , pixel_11_24_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_25_o    , pixel_09_25_o    , pixel_10_25_o    , pixel_11_25_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_26_o    , pixel_09_26_o    , pixel_10_26_o    , pixel_11_26_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_27_o    , pixel_09_27_o    , pixel_10_27_o    , pixel_11_27_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_28_o    , pixel_09_28_o    , pixel_10_28_o    , pixel_11_28_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_29_o    , pixel_09_29_o    , pixel_10_29_o    , pixel_11_29_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_08_30_o    , pixel_09_30_o    , pixel_10_30_o    , pixel_11_30_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_31_o    , pixel_09_31_o    , pixel_10_31_o    , pixel_11_31_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_32_o    , pixel_09_32_o    , pixel_10_32_o    , pixel_11_32_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_33_o    , pixel_09_33_o    , pixel_10_33_o    , pixel_11_33_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_34_o    , pixel_09_34_o    , pixel_10_34_o    , pixel_11_34_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_35_o    , pixel_09_35_o    , pixel_10_35_o    , pixel_11_35_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_36_o    , pixel_09_36_o    , pixel_10_36_o    , pixel_11_36_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_37_o    , pixel_09_37_o    , pixel_10_37_o    , pixel_11_37_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_38_o    , pixel_09_38_o    , pixel_10_38_o    , pixel_11_38_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_39_o    , pixel_09_39_o    , pixel_10_39_o    , pixel_11_39_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_08_40_o    , pixel_09_40_o    , pixel_10_40_o    , pixel_11_40_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_41_o    , pixel_09_41_o    , pixel_10_41_o    , pixel_11_41_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_42_o    , pixel_09_42_o    , pixel_10_42_o    , pixel_11_42_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_43_o    , pixel_09_43_o    , pixel_10_43_o    , pixel_11_43_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_44_o    , pixel_09_44_o    , pixel_10_44_o    , pixel_11_44_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_45_o    , pixel_09_45_o    , pixel_10_45_o    , pixel_11_45_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_46_o    , pixel_09_46_o    , pixel_10_46_o    , pixel_11_46_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_47_o    , pixel_09_47_o    , pixel_10_47_o    , pixel_11_47_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_48_o    , pixel_09_48_o    , pixel_10_48_o    , pixel_11_48_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_49_o    , pixel_09_49_o    , pixel_10_49_o    , pixel_11_49_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_08_50_o    , pixel_09_50_o    , pixel_10_50_o    , pixel_11_50_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_51_o    , pixel_09_51_o    , pixel_10_51_o    , pixel_11_51_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_52_o    , pixel_09_52_o    , pixel_10_52_o    , pixel_11_52_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_53_o    , pixel_09_53_o    , pixel_10_53_o    , pixel_11_53_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_54_o    , pixel_09_54_o    , pixel_10_54_o    , pixel_11_54_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_55_o    , pixel_09_55_o    , pixel_10_55_o    , pixel_11_55_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_56_o    , pixel_09_56_o    , pixel_10_56_o    , pixel_11_56_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_57_o    , pixel_09_57_o    , pixel_10_57_o    , pixel_11_57_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_58_o    , pixel_09_58_o    , pixel_10_58_o    , pixel_11_58_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_59_o    , pixel_09_59_o    , pixel_10_59_o    , pixel_11_59_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_08_60_o    , pixel_09_60_o    , pixel_10_60_o    , pixel_11_60_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_61_o    , pixel_09_61_o    , pixel_10_61_o    , pixel_11_61_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_62_o    , pixel_09_62_o    , pixel_10_62_o    , pixel_11_62_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_08_63_o    , pixel_09_63_o    , pixel_10_63_o    , pixel_11_63_o    ;

  // pixel_12-15_00-63_o
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_00_o    , pixel_13_00_o    , pixel_14_00_o    , pixel_15_00_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_01_o    , pixel_13_01_o    , pixel_14_01_o    , pixel_15_01_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_02_o    , pixel_13_02_o    , pixel_14_02_o    , pixel_15_02_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_03_o    , pixel_13_03_o    , pixel_14_03_o    , pixel_15_03_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_04_o    , pixel_13_04_o    , pixel_14_04_o    , pixel_15_04_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_05_o    , pixel_13_05_o    , pixel_14_05_o    , pixel_15_05_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_06_o    , pixel_13_06_o    , pixel_14_06_o    , pixel_15_06_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_07_o    , pixel_13_07_o    , pixel_14_07_o    , pixel_15_07_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_08_o    , pixel_13_08_o    , pixel_14_08_o    , pixel_15_08_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_09_o    , pixel_13_09_o    , pixel_14_09_o    , pixel_15_09_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_12_10_o    , pixel_13_10_o    , pixel_14_10_o    , pixel_15_10_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_11_o    , pixel_13_11_o    , pixel_14_11_o    , pixel_15_11_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_12_o    , pixel_13_12_o    , pixel_14_12_o    , pixel_15_12_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_13_o    , pixel_13_13_o    , pixel_14_13_o    , pixel_15_13_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_14_o    , pixel_13_14_o    , pixel_14_14_o    , pixel_15_14_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_15_o    , pixel_13_15_o    , pixel_14_15_o    , pixel_15_15_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_16_o    , pixel_13_16_o    , pixel_14_16_o    , pixel_15_16_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_17_o    , pixel_13_17_o    , pixel_14_17_o    , pixel_15_17_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_18_o    , pixel_13_18_o    , pixel_14_18_o    , pixel_15_18_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_19_o    , pixel_13_19_o    , pixel_14_19_o    , pixel_15_19_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_12_20_o    , pixel_13_20_o    , pixel_14_20_o    , pixel_15_20_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_21_o    , pixel_13_21_o    , pixel_14_21_o    , pixel_15_21_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_22_o    , pixel_13_22_o    , pixel_14_22_o    , pixel_15_22_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_23_o    , pixel_13_23_o    , pixel_14_23_o    , pixel_15_23_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_24_o    , pixel_13_24_o    , pixel_14_24_o    , pixel_15_24_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_25_o    , pixel_13_25_o    , pixel_14_25_o    , pixel_15_25_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_26_o    , pixel_13_26_o    , pixel_14_26_o    , pixel_15_26_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_27_o    , pixel_13_27_o    , pixel_14_27_o    , pixel_15_27_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_28_o    , pixel_13_28_o    , pixel_14_28_o    , pixel_15_28_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_29_o    , pixel_13_29_o    , pixel_14_29_o    , pixel_15_29_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_12_30_o    , pixel_13_30_o    , pixel_14_30_o    , pixel_15_30_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_31_o    , pixel_13_31_o    , pixel_14_31_o    , pixel_15_31_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_32_o    , pixel_13_32_o    , pixel_14_32_o    , pixel_15_32_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_33_o    , pixel_13_33_o    , pixel_14_33_o    , pixel_15_33_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_34_o    , pixel_13_34_o    , pixel_14_34_o    , pixel_15_34_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_35_o    , pixel_13_35_o    , pixel_14_35_o    , pixel_15_35_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_36_o    , pixel_13_36_o    , pixel_14_36_o    , pixel_15_36_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_37_o    , pixel_13_37_o    , pixel_14_37_o    , pixel_15_37_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_38_o    , pixel_13_38_o    , pixel_14_38_o    , pixel_15_38_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_39_o    , pixel_13_39_o    , pixel_14_39_o    , pixel_15_39_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_12_40_o    , pixel_13_40_o    , pixel_14_40_o    , pixel_15_40_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_41_o    , pixel_13_41_o    , pixel_14_41_o    , pixel_15_41_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_42_o    , pixel_13_42_o    , pixel_14_42_o    , pixel_15_42_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_43_o    , pixel_13_43_o    , pixel_14_43_o    , pixel_15_43_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_44_o    , pixel_13_44_o    , pixel_14_44_o    , pixel_15_44_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_45_o    , pixel_13_45_o    , pixel_14_45_o    , pixel_15_45_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_46_o    , pixel_13_46_o    , pixel_14_46_o    , pixel_15_46_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_47_o    , pixel_13_47_o    , pixel_14_47_o    , pixel_15_47_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_48_o    , pixel_13_48_o    , pixel_14_48_o    , pixel_15_48_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_49_o    , pixel_13_49_o    , pixel_14_49_o    , pixel_15_49_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_12_50_o    , pixel_13_50_o    , pixel_14_50_o    , pixel_15_50_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_51_o    , pixel_13_51_o    , pixel_14_51_o    , pixel_15_51_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_52_o    , pixel_13_52_o    , pixel_14_52_o    , pixel_15_52_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_53_o    , pixel_13_53_o    , pixel_14_53_o    , pixel_15_53_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_54_o    , pixel_13_54_o    , pixel_14_54_o    , pixel_15_54_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_55_o    , pixel_13_55_o    , pixel_14_55_o    , pixel_15_55_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_56_o    , pixel_13_56_o    , pixel_14_56_o    , pixel_15_56_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_57_o    , pixel_13_57_o    , pixel_14_57_o    , pixel_15_57_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_58_o    , pixel_13_58_o    , pixel_14_58_o    , pixel_15_58_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_59_o    , pixel_13_59_o    , pixel_14_59_o    , pixel_15_59_o    ;

  output [`PIXEL_WIDTH-1    : 0]    pixel_12_60_o    , pixel_13_60_o    , pixel_14_60_o    , pixel_15_60_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_61_o    , pixel_13_61_o    , pixel_14_61_o    , pixel_15_61_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_62_o    , pixel_13_62_o    , pixel_14_62_o    , pixel_15_62_o    ;
  output [`PIXEL_WIDTH-1    : 0]    pixel_12_63_o    , pixel_13_63_o    , pixel_14_63_o    , pixel_15_63_o    ;
*/

//*** WIRE & REG DECLARATION ***************************************************

  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_00_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_01_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_02_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_03_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_04_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_05_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_06_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_07_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_08_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_09_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_10_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_11_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_12_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_13_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_14_r      ;
  reg    [`PIXEL_WIDTH*64-1 : 0]    pixel_15_r      ;


//*** MAIN BODY ****************************************************************

  always @(posedge clk or negedge rstn ) begin
    if( !rstn ) begin
      pixel_00_r <= 'd0 ;
      pixel_01_r <= 'd0 ;
      pixel_02_r <= 'd0 ;
      pixel_03_r <= 'd0 ;
      pixel_04_r <= 'd0 ;
      pixel_05_r <= 'd0 ;
      pixel_06_r <= 'd0 ;
      pixel_07_r <= 'd0 ;
      pixel_08_r <= 'd0 ;
      pixel_09_r <= 'd0 ;
      pixel_10_r <= 'd0 ;
      pixel_11_r <= 'd0 ;
      pixel_12_r <= 'd0 ;
      pixel_13_r <= 'd0 ;
      pixel_14_r <= 'd0 ;
      pixel_15_r <= 'd0 ;
    end
    else if( shift_en_i ) begin
      pixel_15_r <= shift_data_i ;
      pixel_14_r <= pixel_15_r ;
      pixel_13_r <= pixel_14_r ;
      pixel_12_r <= pixel_13_r ;
      pixel_11_r <= pixel_12_r ;
      pixel_10_r <= pixel_11_r ;
      pixel_09_r <= pixel_10_r ;
      pixel_08_r <= pixel_09_r ;
      pixel_07_r <= pixel_08_r ;
      pixel_06_r <= pixel_07_r ;
      pixel_05_r <= pixel_06_r ;
      pixel_04_r <= pixel_05_r ;
      pixel_03_r <= pixel_04_r ;
      pixel_02_r <= pixel_03_r ;
      pixel_01_r <= pixel_02_r ;
      pixel_00_r <= pixel_01_r ;
    end
  end

  assign pixel_00_o = pixel_00_r ;
  assign pixel_01_o = pixel_01_r ;
  assign pixel_02_o = pixel_02_r ;
  assign pixel_03_o = pixel_03_r ;
  assign pixel_04_o = pixel_04_r ;
  assign pixel_05_o = pixel_05_r ;
  assign pixel_06_o = pixel_06_r ;
  assign pixel_07_o = pixel_07_r ;
  assign pixel_08_o = pixel_08_r ;
  assign pixel_09_o = pixel_09_r ;
  assign pixel_10_o = pixel_10_r ;
  assign pixel_11_o = pixel_11_r ;
  assign pixel_12_o = pixel_12_r ;
  assign pixel_13_o = pixel_13_r ;
  assign pixel_14_o = pixel_14_r ;
  assign pixel_15_o = pixel_15_r ;

/*
  assign { pixel_00_00_o ,pixel_00_01_o ,pixel_00_02_o ,pixel_00_03_o ,pixel_00_04_o ,pixel_00_05_o ,pixel_00_06_o ,pixel_00_07_o,
           pixel_00_08_o ,pixel_00_09_o ,pixel_00_10_o ,pixel_00_11_o ,pixel_00_12_o ,pixel_00_13_o ,pixel_00_14_o ,pixel_00_15_o,
           pixel_00_16_o ,pixel_00_17_o ,pixel_00_18_o ,pixel_00_19_o ,pixel_00_20_o ,pixel_00_21_o ,pixel_00_22_o ,pixel_00_23_o,
           pixel_00_24_o ,pixel_00_25_o ,pixel_00_26_o ,pixel_00_27_o ,pixel_00_28_o ,pixel_00_29_o ,pixel_00_30_o ,pixel_00_31_o,
           pixel_00_32_o ,pixel_00_33_o ,pixel_00_34_o ,pixel_00_35_o ,pixel_00_36_o ,pixel_00_37_o ,pixel_00_38_o ,pixel_00_39_o,
           pixel_00_40_o ,pixel_00_41_o ,pixel_00_42_o ,pixel_00_43_o ,pixel_00_44_o ,pixel_00_45_o ,pixel_00_46_o ,pixel_00_47_o,
           pixel_00_48_o ,pixel_00_49_o ,pixel_00_50_o ,pixel_00_51_o ,pixel_00_52_o ,pixel_00_53_o ,pixel_00_54_o ,pixel_00_55_o,
           pixel_00_56_o ,pixel_00_57_o ,pixel_00_58_o ,pixel_00_59_o ,pixel_00_60_o ,pixel_00_61_o ,pixel_00_62_o ,pixel_00_63_o
         } = pixel_00_r ;
         
  assign { pixel_01_00_o ,pixel_01_01_o ,pixel_01_02_o ,pixel_01_03_o ,pixel_01_04_o ,pixel_01_05_o ,pixel_01_06_o ,pixel_01_07_o,
           pixel_01_08_o ,pixel_01_09_o ,pixel_01_10_o ,pixel_01_11_o ,pixel_01_12_o ,pixel_01_13_o ,pixel_01_14_o ,pixel_01_15_o,
           pixel_01_16_o ,pixel_01_17_o ,pixel_01_18_o ,pixel_01_19_o ,pixel_01_20_o ,pixel_01_21_o ,pixel_01_22_o ,pixel_01_23_o,
           pixel_01_24_o ,pixel_01_25_o ,pixel_01_26_o ,pixel_01_27_o ,pixel_01_28_o ,pixel_01_29_o ,pixel_01_30_o ,pixel_01_31_o,
           pixel_01_32_o ,pixel_01_33_o ,pixel_01_34_o ,pixel_01_35_o ,pixel_01_36_o ,pixel_01_37_o ,pixel_01_38_o ,pixel_01_39_o,
           pixel_01_40_o ,pixel_01_41_o ,pixel_01_42_o ,pixel_01_43_o ,pixel_01_44_o ,pixel_01_45_o ,pixel_01_46_o ,pixel_01_47_o,
           pixel_01_48_o ,pixel_01_49_o ,pixel_01_50_o ,pixel_01_51_o ,pixel_01_52_o ,pixel_01_53_o ,pixel_01_54_o ,pixel_01_55_o,
           pixel_01_56_o ,pixel_01_57_o ,pixel_01_58_o ,pixel_01_59_o ,pixel_01_60_o ,pixel_01_61_o ,pixel_01_62_o ,pixel_01_63_o
         } = pixel_01_r ;

  assign { pixel_02_00_o ,pixel_02_01_o ,pixel_02_02_o ,pixel_02_03_o ,pixel_02_04_o ,pixel_02_05_o ,pixel_02_06_o ,pixel_02_07_o,
           pixel_02_08_o ,pixel_02_09_o ,pixel_02_10_o ,pixel_02_11_o ,pixel_02_12_o ,pixel_02_13_o ,pixel_02_14_o ,pixel_02_15_o,
           pixel_02_16_o ,pixel_02_17_o ,pixel_02_18_o ,pixel_02_19_o ,pixel_02_20_o ,pixel_02_21_o ,pixel_02_22_o ,pixel_02_23_o,
           pixel_02_24_o ,pixel_02_25_o ,pixel_02_26_o ,pixel_02_27_o ,pixel_02_28_o ,pixel_02_29_o ,pixel_02_30_o ,pixel_02_31_o,
           pixel_02_32_o ,pixel_02_33_o ,pixel_02_34_o ,pixel_02_35_o ,pixel_02_36_o ,pixel_02_37_o ,pixel_02_38_o ,pixel_02_39_o,
           pixel_02_40_o ,pixel_02_41_o ,pixel_02_42_o ,pixel_02_43_o ,pixel_02_44_o ,pixel_02_45_o ,pixel_02_46_o ,pixel_02_47_o,
           pixel_02_48_o ,pixel_02_49_o ,pixel_02_50_o ,pixel_02_51_o ,pixel_02_52_o ,pixel_02_53_o ,pixel_02_54_o ,pixel_02_55_o,
           pixel_02_56_o ,pixel_02_57_o ,pixel_02_58_o ,pixel_02_59_o ,pixel_02_60_o ,pixel_02_61_o ,pixel_02_62_o ,pixel_02_63_o
         } = pixel_02_r ;

  assign { pixel_03_00_o ,pixel_03_01_o ,pixel_03_02_o ,pixel_03_03_o ,pixel_03_04_o ,pixel_03_05_o ,pixel_03_06_o ,pixel_03_07_o,
           pixel_03_08_o ,pixel_03_09_o ,pixel_03_10_o ,pixel_03_11_o ,pixel_03_12_o ,pixel_03_13_o ,pixel_03_14_o ,pixel_03_15_o,
           pixel_03_16_o ,pixel_03_17_o ,pixel_03_18_o ,pixel_03_19_o ,pixel_03_20_o ,pixel_03_21_o ,pixel_03_22_o ,pixel_03_23_o,
           pixel_03_24_o ,pixel_03_25_o ,pixel_03_26_o ,pixel_03_27_o ,pixel_03_28_o ,pixel_03_29_o ,pixel_03_30_o ,pixel_03_31_o,
           pixel_03_32_o ,pixel_03_33_o ,pixel_03_34_o ,pixel_03_35_o ,pixel_03_36_o ,pixel_03_37_o ,pixel_03_38_o ,pixel_03_39_o,
           pixel_03_40_o ,pixel_03_41_o ,pixel_03_42_o ,pixel_03_43_o ,pixel_03_44_o ,pixel_03_45_o ,pixel_03_46_o ,pixel_03_47_o,
           pixel_03_48_o ,pixel_03_49_o ,pixel_03_50_o ,pixel_03_51_o ,pixel_03_52_o ,pixel_03_53_o ,pixel_03_54_o ,pixel_03_55_o,
           pixel_03_56_o ,pixel_03_57_o ,pixel_03_58_o ,pixel_03_59_o ,pixel_03_60_o ,pixel_03_61_o ,pixel_03_62_o ,pixel_03_63_o
         } = pixel_03_r ;

  assign { pixel_04_00_o ,pixel_04_01_o ,pixel_04_02_o ,pixel_04_03_o ,pixel_04_04_o ,pixel_04_05_o ,pixel_04_06_o ,pixel_04_07_o,
           pixel_04_08_o ,pixel_04_09_o ,pixel_04_10_o ,pixel_04_11_o ,pixel_04_12_o ,pixel_04_13_o ,pixel_04_14_o ,pixel_04_15_o,
           pixel_04_16_o ,pixel_04_17_o ,pixel_04_18_o ,pixel_04_19_o ,pixel_04_20_o ,pixel_04_21_o ,pixel_04_22_o ,pixel_04_23_o,
           pixel_04_24_o ,pixel_04_25_o ,pixel_04_26_o ,pixel_04_27_o ,pixel_04_28_o ,pixel_04_29_o ,pixel_04_30_o ,pixel_04_31_o,
           pixel_04_32_o ,pixel_04_33_o ,pixel_04_34_o ,pixel_04_35_o ,pixel_04_36_o ,pixel_04_37_o ,pixel_04_38_o ,pixel_04_39_o,
           pixel_04_40_o ,pixel_04_41_o ,pixel_04_42_o ,pixel_04_43_o ,pixel_04_44_o ,pixel_04_45_o ,pixel_04_46_o ,pixel_04_47_o,
           pixel_04_48_o ,pixel_04_49_o ,pixel_04_50_o ,pixel_04_51_o ,pixel_04_52_o ,pixel_04_53_o ,pixel_04_54_o ,pixel_04_55_o,
           pixel_04_56_o ,pixel_04_57_o ,pixel_04_58_o ,pixel_04_59_o ,pixel_04_60_o ,pixel_04_61_o ,pixel_04_62_o ,pixel_04_63_o
         } = pixel_04_r ;

  assign { pixel_05_00_o ,pixel_05_01_o ,pixel_05_02_o ,pixel_05_03_o ,pixel_05_04_o ,pixel_05_05_o ,pixel_05_06_o ,pixel_05_07_o,
           pixel_05_08_o ,pixel_05_09_o ,pixel_05_10_o ,pixel_05_11_o ,pixel_05_12_o ,pixel_05_13_o ,pixel_05_14_o ,pixel_05_15_o,
           pixel_05_16_o ,pixel_05_17_o ,pixel_05_18_o ,pixel_05_19_o ,pixel_05_20_o ,pixel_05_21_o ,pixel_05_22_o ,pixel_05_23_o,
           pixel_05_24_o ,pixel_05_25_o ,pixel_05_26_o ,pixel_05_27_o ,pixel_05_28_o ,pixel_05_29_o ,pixel_05_30_o ,pixel_05_31_o,
           pixel_05_32_o ,pixel_05_33_o ,pixel_05_34_o ,pixel_05_35_o ,pixel_05_36_o ,pixel_05_37_o ,pixel_05_38_o ,pixel_05_39_o,
           pixel_05_40_o ,pixel_05_41_o ,pixel_05_42_o ,pixel_05_43_o ,pixel_05_44_o ,pixel_05_45_o ,pixel_05_46_o ,pixel_05_47_o,
           pixel_05_48_o ,pixel_05_49_o ,pixel_05_50_o ,pixel_05_51_o ,pixel_05_52_o ,pixel_05_53_o ,pixel_05_54_o ,pixel_05_55_o,
           pixel_05_56_o ,pixel_05_57_o ,pixel_05_58_o ,pixel_05_59_o ,pixel_05_60_o ,pixel_05_61_o ,pixel_05_62_o ,pixel_05_63_o
         } = pixel_05_r ;

  assign { pixel_06_00_o ,pixel_06_01_o ,pixel_06_02_o ,pixel_06_03_o ,pixel_06_04_o ,pixel_06_05_o ,pixel_06_06_o ,pixel_06_07_o,
           pixel_06_08_o ,pixel_06_09_o ,pixel_06_10_o ,pixel_06_11_o ,pixel_06_12_o ,pixel_06_13_o ,pixel_06_14_o ,pixel_06_15_o,
           pixel_06_16_o ,pixel_06_17_o ,pixel_06_18_o ,pixel_06_19_o ,pixel_06_20_o ,pixel_06_21_o ,pixel_06_22_o ,pixel_06_23_o,
           pixel_06_24_o ,pixel_06_25_o ,pixel_06_26_o ,pixel_06_27_o ,pixel_06_28_o ,pixel_06_29_o ,pixel_06_30_o ,pixel_06_31_o,
           pixel_06_32_o ,pixel_06_33_o ,pixel_06_34_o ,pixel_06_35_o ,pixel_06_36_o ,pixel_06_37_o ,pixel_06_38_o ,pixel_06_39_o,
           pixel_06_40_o ,pixel_06_41_o ,pixel_06_42_o ,pixel_06_43_o ,pixel_06_44_o ,pixel_06_45_o ,pixel_06_46_o ,pixel_06_47_o,
           pixel_06_48_o ,pixel_06_49_o ,pixel_06_50_o ,pixel_06_51_o ,pixel_06_52_o ,pixel_06_53_o ,pixel_06_54_o ,pixel_06_55_o,
           pixel_06_56_o ,pixel_06_57_o ,pixel_06_58_o ,pixel_06_59_o ,pixel_06_60_o ,pixel_06_61_o ,pixel_06_62_o ,pixel_06_63_o
         } = pixel_06_r ;

  assign { pixel_07_00_o ,pixel_07_01_o ,pixel_07_02_o ,pixel_07_03_o ,pixel_07_04_o ,pixel_07_05_o ,pixel_07_06_o ,pixel_07_07_o,
           pixel_07_08_o ,pixel_07_09_o ,pixel_07_10_o ,pixel_07_11_o ,pixel_07_12_o ,pixel_07_13_o ,pixel_07_14_o ,pixel_07_15_o,
           pixel_07_16_o ,pixel_07_17_o ,pixel_07_18_o ,pixel_07_19_o ,pixel_07_20_o ,pixel_07_21_o ,pixel_07_22_o ,pixel_07_23_o,
           pixel_07_24_o ,pixel_07_25_o ,pixel_07_26_o ,pixel_07_27_o ,pixel_07_28_o ,pixel_07_29_o ,pixel_07_30_o ,pixel_07_31_o,
           pixel_07_32_o ,pixel_07_33_o ,pixel_07_34_o ,pixel_07_35_o ,pixel_07_36_o ,pixel_07_37_o ,pixel_07_38_o ,pixel_07_39_o,
           pixel_07_40_o ,pixel_07_41_o ,pixel_07_42_o ,pixel_07_43_o ,pixel_07_44_o ,pixel_07_45_o ,pixel_07_46_o ,pixel_07_47_o,
           pixel_07_48_o ,pixel_07_49_o ,pixel_07_50_o ,pixel_07_51_o ,pixel_07_52_o ,pixel_07_53_o ,pixel_07_54_o ,pixel_07_55_o,
           pixel_07_56_o ,pixel_07_57_o ,pixel_07_58_o ,pixel_07_59_o ,pixel_07_60_o ,pixel_07_61_o ,pixel_07_62_o ,pixel_07_63_o
         } = pixel_07_r ;

  assign { pixel_08_00_o ,pixel_08_01_o ,pixel_08_02_o ,pixel_08_03_o ,pixel_08_04_o ,pixel_08_05_o ,pixel_08_06_o ,pixel_08_07_o,
           pixel_08_08_o ,pixel_08_09_o ,pixel_08_10_o ,pixel_08_11_o ,pixel_08_12_o ,pixel_08_13_o ,pixel_08_14_o ,pixel_08_15_o,
           pixel_08_16_o ,pixel_08_17_o ,pixel_08_18_o ,pixel_08_19_o ,pixel_08_20_o ,pixel_08_21_o ,pixel_08_22_o ,pixel_08_23_o,
           pixel_08_24_o ,pixel_08_25_o ,pixel_08_26_o ,pixel_08_27_o ,pixel_08_28_o ,pixel_08_29_o ,pixel_08_30_o ,pixel_08_31_o,
           pixel_08_32_o ,pixel_08_33_o ,pixel_08_34_o ,pixel_08_35_o ,pixel_08_36_o ,pixel_08_37_o ,pixel_08_38_o ,pixel_08_39_o,
           pixel_08_40_o ,pixel_08_41_o ,pixel_08_42_o ,pixel_08_43_o ,pixel_08_44_o ,pixel_08_45_o ,pixel_08_46_o ,pixel_08_47_o,
           pixel_08_48_o ,pixel_08_49_o ,pixel_08_50_o ,pixel_08_51_o ,pixel_08_52_o ,pixel_08_53_o ,pixel_08_54_o ,pixel_08_55_o,
           pixel_08_56_o ,pixel_08_57_o ,pixel_08_58_o ,pixel_08_59_o ,pixel_08_60_o ,pixel_08_61_o ,pixel_08_62_o ,pixel_08_63_o
         } = pixel_08_r ;

  assign { pixel_09_00_o ,pixel_09_01_o ,pixel_09_02_o ,pixel_09_03_o ,pixel_09_04_o ,pixel_09_05_o ,pixel_09_06_o ,pixel_09_07_o,
           pixel_09_08_o ,pixel_09_09_o ,pixel_09_10_o ,pixel_09_11_o ,pixel_09_12_o ,pixel_09_13_o ,pixel_09_14_o ,pixel_09_15_o,
           pixel_09_16_o ,pixel_09_17_o ,pixel_09_18_o ,pixel_09_19_o ,pixel_09_20_o ,pixel_09_21_o ,pixel_09_22_o ,pixel_09_23_o,
           pixel_09_24_o ,pixel_09_25_o ,pixel_09_26_o ,pixel_09_27_o ,pixel_09_28_o ,pixel_09_29_o ,pixel_09_30_o ,pixel_09_31_o,
           pixel_09_32_o ,pixel_09_33_o ,pixel_09_34_o ,pixel_09_35_o ,pixel_09_36_o ,pixel_09_37_o ,pixel_09_38_o ,pixel_09_39_o,
           pixel_09_40_o ,pixel_09_41_o ,pixel_09_42_o ,pixel_09_43_o ,pixel_09_44_o ,pixel_09_45_o ,pixel_09_46_o ,pixel_09_47_o,
           pixel_09_48_o ,pixel_09_49_o ,pixel_09_50_o ,pixel_09_51_o ,pixel_09_52_o ,pixel_09_53_o ,pixel_09_54_o ,pixel_09_55_o,
           pixel_09_56_o ,pixel_09_57_o ,pixel_09_58_o ,pixel_09_59_o ,pixel_09_60_o ,pixel_09_61_o ,pixel_09_62_o ,pixel_09_63_o
         } = pixel_09_r ;

  assign { pixel_10_00_o ,pixel_10_01_o ,pixel_10_02_o ,pixel_10_03_o ,pixel_10_04_o ,pixel_10_05_o ,pixel_10_06_o ,pixel_10_07_o,
           pixel_10_08_o ,pixel_10_09_o ,pixel_10_10_o ,pixel_10_11_o ,pixel_10_12_o ,pixel_10_13_o ,pixel_10_14_o ,pixel_10_15_o,
           pixel_10_16_o ,pixel_10_17_o ,pixel_10_18_o ,pixel_10_19_o ,pixel_10_20_o ,pixel_10_21_o ,pixel_10_22_o ,pixel_10_23_o,
           pixel_10_24_o ,pixel_10_25_o ,pixel_10_26_o ,pixel_10_27_o ,pixel_10_28_o ,pixel_10_29_o ,pixel_10_30_o ,pixel_10_31_o,
           pixel_10_32_o ,pixel_10_33_o ,pixel_10_34_o ,pixel_10_35_o ,pixel_10_36_o ,pixel_10_37_o ,pixel_10_38_o ,pixel_10_39_o,
           pixel_10_40_o ,pixel_10_41_o ,pixel_10_42_o ,pixel_10_43_o ,pixel_10_44_o ,pixel_10_45_o ,pixel_10_46_o ,pixel_10_47_o,
           pixel_10_48_o ,pixel_10_49_o ,pixel_10_50_o ,pixel_10_51_o ,pixel_10_52_o ,pixel_10_53_o ,pixel_10_54_o ,pixel_10_55_o,
           pixel_10_56_o ,pixel_10_57_o ,pixel_10_58_o ,pixel_10_59_o ,pixel_10_60_o ,pixel_10_61_o ,pixel_10_62_o ,pixel_10_63_o
         } = pixel_10_r ;

  assign { pixel_11_00_o ,pixel_11_01_o ,pixel_11_02_o ,pixel_11_03_o ,pixel_11_04_o ,pixel_11_05_o ,pixel_11_06_o ,pixel_11_07_o,
           pixel_11_08_o ,pixel_11_09_o ,pixel_11_10_o ,pixel_11_11_o ,pixel_11_12_o ,pixel_11_13_o ,pixel_11_14_o ,pixel_11_15_o,
           pixel_11_16_o ,pixel_11_17_o ,pixel_11_18_o ,pixel_11_19_o ,pixel_11_20_o ,pixel_11_21_o ,pixel_11_22_o ,pixel_11_23_o,
           pixel_11_24_o ,pixel_11_25_o ,pixel_11_26_o ,pixel_11_27_o ,pixel_11_28_o ,pixel_11_29_o ,pixel_11_30_o ,pixel_11_31_o,
           pixel_11_32_o ,pixel_11_33_o ,pixel_11_34_o ,pixel_11_35_o ,pixel_11_36_o ,pixel_11_37_o ,pixel_11_38_o ,pixel_11_39_o,
           pixel_11_40_o ,pixel_11_41_o ,pixel_11_42_o ,pixel_11_43_o ,pixel_11_44_o ,pixel_11_45_o ,pixel_11_46_o ,pixel_11_47_o,
           pixel_11_48_o ,pixel_11_49_o ,pixel_11_50_o ,pixel_11_51_o ,pixel_11_52_o ,pixel_11_53_o ,pixel_11_54_o ,pixel_11_55_o,
           pixel_11_56_o ,pixel_11_57_o ,pixel_11_58_o ,pixel_11_59_o ,pixel_11_60_o ,pixel_11_61_o ,pixel_11_62_o ,pixel_11_63_o
         } = pixel_11_r ;

  assign { pixel_12_00_o ,pixel_12_01_o ,pixel_12_02_o ,pixel_12_03_o ,pixel_12_04_o ,pixel_12_05_o ,pixel_12_06_o ,pixel_12_07_o,
           pixel_12_08_o ,pixel_12_09_o ,pixel_12_10_o ,pixel_12_11_o ,pixel_12_12_o ,pixel_12_13_o ,pixel_12_14_o ,pixel_12_15_o,
           pixel_12_16_o ,pixel_12_17_o ,pixel_12_18_o ,pixel_12_19_o ,pixel_12_20_o ,pixel_12_21_o ,pixel_12_22_o ,pixel_12_23_o,
           pixel_12_24_o ,pixel_12_25_o ,pixel_12_26_o ,pixel_12_27_o ,pixel_12_28_o ,pixel_12_29_o ,pixel_12_30_o ,pixel_12_31_o,
           pixel_12_32_o ,pixel_12_33_o ,pixel_12_34_o ,pixel_12_35_o ,pixel_12_36_o ,pixel_12_37_o ,pixel_12_38_o ,pixel_12_39_o,
           pixel_12_40_o ,pixel_12_41_o ,pixel_12_42_o ,pixel_12_43_o ,pixel_12_44_o ,pixel_12_45_o ,pixel_12_46_o ,pixel_12_47_o,
           pixel_12_48_o ,pixel_12_49_o ,pixel_12_50_o ,pixel_12_51_o ,pixel_12_52_o ,pixel_12_53_o ,pixel_12_54_o ,pixel_12_55_o,
           pixel_12_56_o ,pixel_12_57_o ,pixel_12_58_o ,pixel_12_59_o ,pixel_12_60_o ,pixel_12_61_o ,pixel_12_62_o ,pixel_12_63_o
         } = pixel_12_r ;

  assign { pixel_13_00_o ,pixel_13_01_o ,pixel_13_02_o ,pixel_13_03_o ,pixel_13_04_o ,pixel_13_05_o ,pixel_13_06_o ,pixel_13_07_o,
           pixel_13_08_o ,pixel_13_09_o ,pixel_13_10_o ,pixel_13_11_o ,pixel_13_12_o ,pixel_13_13_o ,pixel_13_14_o ,pixel_13_15_o,
           pixel_13_16_o ,pixel_13_17_o ,pixel_13_18_o ,pixel_13_19_o ,pixel_13_20_o ,pixel_13_21_o ,pixel_13_22_o ,pixel_13_23_o,
           pixel_13_24_o ,pixel_13_25_o ,pixel_13_26_o ,pixel_13_27_o ,pixel_13_28_o ,pixel_13_29_o ,pixel_13_30_o ,pixel_13_31_o,
           pixel_13_32_o ,pixel_13_33_o ,pixel_13_34_o ,pixel_13_35_o ,pixel_13_36_o ,pixel_13_37_o ,pixel_13_38_o ,pixel_13_39_o,
           pixel_13_40_o ,pixel_13_41_o ,pixel_13_42_o ,pixel_13_43_o ,pixel_13_44_o ,pixel_13_45_o ,pixel_13_46_o ,pixel_13_47_o,
           pixel_13_48_o ,pixel_13_49_o ,pixel_13_50_o ,pixel_13_51_o ,pixel_13_52_o ,pixel_13_53_o ,pixel_13_54_o ,pixel_13_55_o,
           pixel_13_56_o ,pixel_13_57_o ,pixel_13_58_o ,pixel_13_59_o ,pixel_13_60_o ,pixel_13_61_o ,pixel_13_62_o ,pixel_13_63_o
         } = pixel_13_r ;

  assign { pixel_14_00_o ,pixel_14_01_o ,pixel_14_02_o ,pixel_14_03_o ,pixel_14_04_o ,pixel_14_05_o ,pixel_14_06_o ,pixel_14_07_o,
           pixel_14_08_o ,pixel_14_09_o ,pixel_14_10_o ,pixel_14_11_o ,pixel_14_12_o ,pixel_14_13_o ,pixel_14_14_o ,pixel_14_15_o,
           pixel_14_16_o ,pixel_14_17_o ,pixel_14_18_o ,pixel_14_19_o ,pixel_14_20_o ,pixel_14_21_o ,pixel_14_22_o ,pixel_14_23_o,
           pixel_14_24_o ,pixel_14_25_o ,pixel_14_26_o ,pixel_14_27_o ,pixel_14_28_o ,pixel_14_29_o ,pixel_14_30_o ,pixel_14_31_o,
           pixel_14_32_o ,pixel_14_33_o ,pixel_14_34_o ,pixel_14_35_o ,pixel_14_36_o ,pixel_14_37_o ,pixel_14_38_o ,pixel_14_39_o,
           pixel_14_40_o ,pixel_14_41_o ,pixel_14_42_o ,pixel_14_43_o ,pixel_14_44_o ,pixel_14_45_o ,pixel_14_46_o ,pixel_14_47_o,
           pixel_14_48_o ,pixel_14_49_o ,pixel_14_50_o ,pixel_14_51_o ,pixel_14_52_o ,pixel_14_53_o ,pixel_14_54_o ,pixel_14_55_o,
           pixel_14_56_o ,pixel_14_57_o ,pixel_14_58_o ,pixel_14_59_o ,pixel_14_60_o ,pixel_14_61_o ,pixel_14_62_o ,pixel_14_63_o
         } = pixel_14_r ;

  assign { pixel_15_00_o ,pixel_15_01_o ,pixel_15_02_o ,pixel_15_03_o ,pixel_15_04_o ,pixel_15_05_o ,pixel_15_06_o ,pixel_15_07_o,
           pixel_15_08_o ,pixel_15_09_o ,pixel_15_10_o ,pixel_15_11_o ,pixel_15_12_o ,pixel_15_13_o ,pixel_15_14_o ,pixel_15_15_o,
           pixel_15_16_o ,pixel_15_17_o ,pixel_15_18_o ,pixel_15_19_o ,pixel_15_20_o ,pixel_15_21_o ,pixel_15_22_o ,pixel_15_23_o,
           pixel_15_24_o ,pixel_15_25_o ,pixel_15_26_o ,pixel_15_27_o ,pixel_15_28_o ,pixel_15_29_o ,pixel_15_30_o ,pixel_15_31_o,
           pixel_15_32_o ,pixel_15_33_o ,pixel_15_34_o ,pixel_15_35_o ,pixel_15_36_o ,pixel_15_37_o ,pixel_15_38_o ,pixel_15_39_o,
           pixel_15_40_o ,pixel_15_41_o ,pixel_15_42_o ,pixel_15_43_o ,pixel_15_44_o ,pixel_15_45_o ,pixel_15_46_o ,pixel_15_47_o,
           pixel_15_48_o ,pixel_15_49_o ,pixel_15_50_o ,pixel_15_51_o ,pixel_15_52_o ,pixel_15_53_o ,pixel_15_54_o ,pixel_15_55_o,
           pixel_15_56_o ,pixel_15_57_o ,pixel_15_58_o ,pixel_15_59_o ,pixel_15_60_o ,pixel_15_61_o ,pixel_15_62_o ,pixel_15_63_o
         } = pixel_15_r ;
*/

//*** DEBUG ********************************************************************


endmodule